`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AGH
// Engineer: Aleksandra Roman, Karolina Brodziak
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_you_win_font
// Project Name: Entliczek pentliczek
// Target Devices: 
// Tool Versions: 
// Description: Du�a czcionka dla napisu YOU WIN
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Wzorowano na czcionce Arcade Classic
//////////////////////////////////////////////////////////////////////////////////


module arcade_you_win_font(
    input  wire        clk,
    input  wire [15:0] addr,            
    output reg  [63:0] char_line_pixels 
);

    // signal declaration
    reg [63:0] data;

// body
always @(posedge clk)
    char_line_pixels <= data;

always @* begin
    case (addr)
        //code x00
        16'h0000: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0001: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0002: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0003: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0004: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0005: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0006: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0007: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0008: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0009: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0010: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0011: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0012: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0013: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0014: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0015: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0016: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0017: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0018: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0019: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0020: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0021: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0022: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0023: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0024: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0025: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0026: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0027: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0028: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0029: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0030: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0031: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0032: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0033: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0034: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0035: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0036: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0037: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0038: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0039: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x4F
        16'h4f00: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f01: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f02: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f03: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f04: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f05: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f06: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f07: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h4f08: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f09: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f10: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f11: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f12: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f13: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f14: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f15: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f16: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f17: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f18: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f19: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f20: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f21: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f22: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f23: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f24: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f25: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f26: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f27: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f28: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f29: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f30: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f31: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f32: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f33: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f34: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f35: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f36: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f37: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h4f38: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f39: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 

        //code x49
        16'h4900: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4901: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4902: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000;  
        16'h4903: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4904: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4905: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4906: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4907: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        
        16'h4908: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4909: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h490a: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h490b: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h490c: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;   
        16'h490d: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h490e: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h490f: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h4910: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4911: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4912: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4913: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4914: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4915: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4916: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;   
        16'h4917: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h4918: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4919: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491a: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491b: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491c: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491d: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491e: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h491f: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h4920: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;   
        16'h4921: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4922: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4923: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4924: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4925: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4926: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4927: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;
        
        16'h4928: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h4929: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h492a: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h492b: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h492c: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h492d: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h492e: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h492f: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h4930: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4931: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4932: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4933: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4934: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000;   
        16'h4935: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4936: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4937: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        
        16'h4938: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4939: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h493a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h493b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h493c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h493d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h493e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;  
        16'h493f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x4e
        16'h4e00: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e01: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e02: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e03: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e04: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e05: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e06: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e07: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4e08: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000;
        16'h4e09: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0a: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0b: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0c: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0d: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0e: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4e0f: data = 64'b11111111_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4e10: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e11: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e12: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e13: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e14: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e15: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e16: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        16'h4e17: data = 64'b11111111_11111111_11111111_11111111_00000000_11111111_11111111_00000000; 
        
        16'h4e18: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e19: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1a: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1b: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1c: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1d: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1e: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4e1f: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        
        16'h4e20: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e21: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e22: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e23: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e24: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e25: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e26: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        16'h4e27: data = 64'b11111111_11111111_00000000_11111111_11111111_11111111_11111111_00000000; 
        
        16'h4e28: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;  
        16'h4e29: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;   
        16'h4e2a: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;  
        16'h4e2b: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;  
        16'h4e2c: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h4e2d: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;   
        16'h4e2e: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h4e2f: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        
        16'h4e30: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e31: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h4e32: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e33: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e34: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e35: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4e36: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4e37: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4e38: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4e39: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4e3a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4e3b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4e3c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4e3d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4e3e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4e3f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x55
        16'h5500: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5501: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5502: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5503: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5504: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5505: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5506: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5507: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5508: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5509: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h550f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5510: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5511: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5512: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5513: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5514: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5515: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5516: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5517: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5518: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5519: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h551f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5520: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5521: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5522: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5523: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5524: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5525: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5526: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5527: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5528: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5529: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h552f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5530: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5531: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5532: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5533: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5534: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5535: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5536: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5537: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h5538: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h5539: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h553f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x57
        16'h5700: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5701: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5702: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5703: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5704: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5705: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5706: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5707: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5708: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5709: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h570f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5710: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5711: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5712: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5713: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5714: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5715: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5716: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5717: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5718: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h5719: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571a: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571b: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571c: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571d: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571e: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        16'h571f: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000; 
        
        16'h5720: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5721: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5722: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5723: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5724: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5725: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5726: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h5727: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        
        16'h5728: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;  
        16'h5729: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;   
        16'h572a: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;  
        16'h572b: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;  
        16'h572c: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000; 
        16'h572d: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;   
        16'h572e: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000; 
        16'h572f: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000; 
        
        16'h5730: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5731: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h5732: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5733: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5734: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5735: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5736: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5737: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5738: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h5739: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h573a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h573b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h573c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h573d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h573e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h573f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x59
        16'h5900: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5901: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000;  
        16'h5902: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5903: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5904: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5905: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5906: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5907: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
       
        16'h5908: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5909: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590a: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590b: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590c: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590d: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590e: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h590f: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5910: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5911: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5912: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5913: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5914: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5915: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5916: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h5917: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5918: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5919: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h591a: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h591b: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h591c: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000;  
        16'h591d: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h591e: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h591f: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000;  
        
        16'h5920: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h5921: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5922: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5923: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5924: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5925: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5926: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5927: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h5928: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5929: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h592a: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h592b: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h592c: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h592d: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h592e: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h592f: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h5930: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5931: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;
        16'h5932: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5933: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5934: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000;  
        16'h5935: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5936: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        16'h5937: data = 64'b00000000_00000000_00000000_11111111_11111111_00000000_00000000_00000000; 
        
        16'h5938: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h5939: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h593a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h593b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h593c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h593d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h593e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;  
        16'h593f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        default: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
    endcase
end

endmodule