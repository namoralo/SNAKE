`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_big_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arcade_small_font(
        input  wire        clk,
        input  wire [15:0] addr,            // {char_code[6:0], char_line[3:0]}
        output reg  [39:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [39:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @* begin
        case (addr)
        //code x00
                16'h0000: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0001: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0002: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0003: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0004: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
                 
                16'h0005: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0006: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0007: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0008: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0009: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                
                16'h000a: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h000b: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h000c: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h000d: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h000e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                
                16'h000f: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0010: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0011: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0012: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0013: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
              
                16'h0014: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0015: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0016: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0017: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0018: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
                 
                16'h0019: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h001a: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h001b: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h001c: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h001d: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
       
                16'h001e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h001f: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0020: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0021: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0022: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                
                16'h0023: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0024: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0025: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0026: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                16'h0027: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
                

                    //code x47
        16'h4700: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
        16'h4701: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
        16'h4702: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
        16'h4703: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
        16'h4704: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;
          
        16'h4705: data = 40'b00000_11111_11111_00000_00000_00000_00000_00000;
        16'h4706: data = 40'b00000_11111_11111_00000_00000_00000_00000_00000; 
        16'h4707: data = 40'b00000_11111_11111_00000_00000_00000_00000_00000; 
        16'h4708: data = 40'b00000_11111_11111_00000_00000_00000_00000_00000; 
        16'h4709: data = 40'b00000_11111_11111_00000_00000_00000_00000_00000; 
        
        16'h470a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
        16'h470b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
        16'h470c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
        16'h470d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
        16'h470e: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;
         
        16'h470f: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
        16'h4710: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
        16'h4711: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
        16'h4712: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
        16'h4713: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
       
        16'h4714: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
        16'h4715: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
        16'h4716: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
        16'h4717: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
        16'h4718: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
        
        16'h4719: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
        16'h471a: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
        16'h471b: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
        16'h471c: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
        16'h471d: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 

        16'h471e: data = 40'b00000_00000_11111_11111_11111_11111_11111_00000; 
        16'h471f: data = 40'b00000_00000_11111_11111_11111_11111_11111_00000; 
        16'h4720: data = 40'b00000_00000_11111_11111_11111_11111_11111_00000; 
        16'h4721: data = 40'b00000_00000_11111_11111_11111_11111_11111_00000; 
        16'h4722: data = 40'b00000_00000_11111_11111_11111_11111_11111_00000;
         
        16'h4723: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        16'h4724: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        16'h4725: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        16'h4726: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        16'h4727: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        
        default: data = 40'b0;
        
          
        endcase
end
endmodule

