`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_big_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arcade_big_font(
        input  wire        clk,
        input  wire [15:0] addr,            // {char_code[6:0], char_line[3:0]}
        output reg  [79:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [79:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @* begin
        case (addr)
        //code x00
                16'h0000: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0001: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0002: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0003: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0004: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0005: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0006: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0007: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0008: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0009: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h000a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0010: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0011: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0012: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0013: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              
                16'h0014: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0015: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0016: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0017: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0018: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0019: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
       
                16'h001e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0020: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0021: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0022: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0023: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0024: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0025: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0026: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0027: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h0028: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0029: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0030: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0031: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        
                16'h0032: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0033: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0034: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0035: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0036: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0037: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0038: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0039: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h003c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0040: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0041: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0042: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0043: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0044: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0045: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                
                16'h0046: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0047: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0048: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0049: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                

                    //code x47
        16'h4700: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4701: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4702: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4703: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4704: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4705: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4706: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4707: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4708: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4709: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        
        16'h470a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470c: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470d: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470e: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470f: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4710: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4711: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4712: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4713: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
       
        16'h4714: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4715: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4716: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4717: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4718: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4719: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 

        16'h471e: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h471f: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4720: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4721: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4722: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4723: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4724: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4725: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4726: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4727: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        
        16'h4728: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4729: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4730: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4731: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 

        16'h4732: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4733: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4734: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4735: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4736: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4737: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4738: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4739: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h473a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h473b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
       
        16'h473c: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473d: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473e: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473f: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4740: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4741: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4742: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4743: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4744: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4745: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        
        16'h4746: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4747: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4748: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4749: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        
        default: data = 80'b0;  
        endcase
end
endmodule

