`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_big_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arcade_game_over_font(
        input  wire        clk,
        input  wire [15:0] addr,            
        output reg  [79:0]  char_line_pixels 
    );

    // signal declaration
    reg [79:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
        //code x00
               16'h0000: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0001: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0002: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0003: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0004: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0005: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0006: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0007: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0008: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0009: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h000a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0010: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0011: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0012: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0013: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              
                16'h0014: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0015: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0016: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0017: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0018: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0019: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
       
                16'h001e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0020: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0021: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0022: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0023: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0024: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0025: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0026: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0027: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h0028: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0029: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0030: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0031: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        
                16'h0032: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0033: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0034: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0035: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0036: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0037: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0038: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0039: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h003c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0040: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0041: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0042: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0043: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0044: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0045: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                
                16'h0046: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0047: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0048: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0049: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;

               //code x41
      16'h4100: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4101: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4102: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4103: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4104: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4105: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4106: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4107: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4108: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
      16'h4109: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;

      16'h410a: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000;
      16'h410b: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h410c: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h410d: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h410e: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h410f: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h4110: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h4111: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h4112: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      16'h4113: data = 80'b0000000000_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000_0000000000; 
      
      16'h4114: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4115: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4116: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4117: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4118: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4119: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h411a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h411b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h411c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h411d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     
      16'h411e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h411f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4120: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4121: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4122: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4123: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4124: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4125: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4126: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4127: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
      
      16'h4128: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
      16'h4129: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412a: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412b: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412c: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412d: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h412f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h4130: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      16'h4131: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
      
      16'h4132: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4133: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4134: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4135: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4136: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4137: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4138: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4139: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h413a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h413b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      
      16'h413c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h413d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h413e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h413f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4140: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4141: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4142: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4143: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4144: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      16'h4145: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
      
      16'h4146: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h4147: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h4148: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h4149: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
      16'h414f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
             
             //code x45
                        16'h4500: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4501: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4502: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4503: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4504: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4505: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4506: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4507: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4508: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4509: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                 
                        16'h450a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h450b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h450c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h450d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h450e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h450f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4510: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4511: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4512: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4513: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                      
                        16'h4514: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4515: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4516: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4517: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4518: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4519: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h451a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h451b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h451c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h451d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        
                        16'h451e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                        16'h451f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        16'h4520: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        16'h4521: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        16'h4522: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                        16'h4523: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                        16'h4524: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        16'h4525: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        16'h4526: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                        16'h4527: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
                        
                        16'h4528: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4529: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;  
                        16'h452a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h452b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h452c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h452d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;  
                        16'h452e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h452f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;  
                        16'h4530: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4531: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                      
                        16'h4532: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4533: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4534: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4535: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4536: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4537: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4538: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
                        16'h4539: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h453a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h453b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        
                        16'h453c: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h453d: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h453e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h453f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                        16'h4540: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h4541: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h4542: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h4543: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h4544: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                        16'h4545: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
                         
                        16'h4546: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4547: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4548: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h4549: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                        16'h454f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;      
                

                    //code x47
        16'h4700: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4701: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4702: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4703: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4704: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4705: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4706: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4707: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4708: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h4709: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        
        16'h470a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470c: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470d: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470e: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h470f: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4710: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4711: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4712: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4713: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000; 
       
        16'h4714: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4715: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4716: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4717: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4718: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4719: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h471d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 

        16'h471e: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h471f: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4720: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4721: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4722: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4723: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4724: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4725: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4726: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        16'h4727: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
        
        16'h4728: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4729: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h472f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4730: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4731: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 

        16'h4732: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4733: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4734: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4735: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4736: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4737: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4738: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h4739: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h473a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h473b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
       
        16'h473c: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473d: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473e: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h473f: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4740: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4741: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4742: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4743: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4744: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        16'h4745: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
        
        16'h4746: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4747: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4748: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h4749: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h474f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
      
        
        
                            //code x4D
              16'h4d00: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d01: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d02: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d03: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d04: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d05: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d06: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d07: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d08: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d09: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                      
              16'h4d0a: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000; 
              16'h4d0b: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d0c: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d0d: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d0e: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d0f: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d10: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d11: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d12: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              16'h4d13: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
              
              16'h4d14: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d15: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d16: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d17: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d18: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d19: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d1a: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d1b: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d1c: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d1d: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
      
              16'h4d1e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d1f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d20: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d21: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d22: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d23: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d24: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d25: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d26: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              16'h4d27: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;
              
              16'h4d28: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d29: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2a: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2b: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2c: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2d: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2e: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d2f: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d30: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
              16'h4d31: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
      
              16'h4d32: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d33: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d34: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d35: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d36: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d37: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d38: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d39: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d3a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d3b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
             
              16'h4d3c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d3d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d3e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d3f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d40: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d41: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d42: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d43: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
              16'h4d44: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              16'h4d45: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              
              16'h4d46: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d47: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d48: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d49: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              16'h4d4f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;  
           
                   //code x4F
     16'h4f00: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f01: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f02: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f03: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f04: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f05: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f06: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f07: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f08: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f09: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     
     16'h4f0a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f10: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f11: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f12: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f13: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
    
     16'h4f14: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f15: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f16: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f17: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f18: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f19: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     
     16'h4f1e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f20: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f21: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f22: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f23: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f24: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f25: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f26: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f27: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     
     16'h4f28: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f29: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f30: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f31: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 

     16'h4f32: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f33: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f34: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f35: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f36: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f37: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f38: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f39: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f3a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f3b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
    
     16'h4f3c: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3d: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3e: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3f: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f40: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f41: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f42: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f43: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f44: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f45: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     
     16'h4f46: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f47: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f48: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f49: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;


                //code x52
                  16'h5200: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5201: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5202: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5203: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5204: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5205: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5206: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5207: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5208: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                  16'h5209: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
           
                  16'h520a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h520b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h520c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h520d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h520e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h520f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5210: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5211: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_11111111110000000000;
                  16'h5212: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5213: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                
                  16'h5214: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5215: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5216: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5217: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5218: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5219: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h521a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h521b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h521c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h521d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                
                  16'h521e: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h521f: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5220: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5221: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5222: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5223: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5224: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5225: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5226: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  16'h5227: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                  
                  16'h5228: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h5229: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;   
                  16'h522a: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h522b: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h522c: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h522d: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;  
                  16'h522e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h522f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;   
                  16'h5230: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                  16'h5231: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
                
                  16'h5232: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h5233: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h5234: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h5235: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h5236: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h5237: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000;
                  16'h5238: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000;
                  16'h5239: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h523a: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  16'h523b: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000; 
                  
                  16'h523c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h523d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h523e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h523f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                  16'h5240: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5241: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5242: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5243: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5244: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                  16'h5245: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                   
                  16'h5246: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h5247: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h5248: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h5249: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                  16'h524f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;      
                       
 //code x56
         16'h5600: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5601: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
         16'h5602: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
         16'h5603: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
         16'h5604: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5605: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5606: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5607: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5608: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
         16'h5609: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
       
         16'h560a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h560b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h560c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h560d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h560e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h560f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5610: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5611: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5612: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5613: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
        
         16'h5614: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5615: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5616: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5617: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5618: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5619: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h561a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h561b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h561c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h561d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         
         16'h561e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h561f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5620: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5621: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5622: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5623: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5624: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5625: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5626: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         16'h5627: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
         
         16'h5628: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h5629: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000;  
         16'h562a: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h562b: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h562c: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h562d: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000;  
         16'h562e: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h562f: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h5630: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
         16'h5631: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
    
         16'h5632: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h5633: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
         16'h5634: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h5635: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
         16'h5636: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h5637: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h5638: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
         16'h5639: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h563a: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000; 
         16'h563b: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000;
        
         16'h563c: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h563d: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h563e: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h563f: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h5640: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000;  
         16'h5641: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h5642: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h5643: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h5644: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000; 
         16'h5645: data = 80'b0000000000_0000000000_0000000000_1111111111_0000000000_0000000000_0000000000_0000000000;  
         
         16'h5646: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h5647: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h5648: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h5649: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
         16'h564f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;

 	default: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        endcase

endmodule

