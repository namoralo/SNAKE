`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: AGH
// Engineer: Aleksandra Roman, Karolina Brodziak
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_game_over_font
// Project Name: Entliczek pentliczek
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Wzorowano na czcionce Arcade Classic
//////////////////////////////////////////////////////////////////////////////////


module arcade_game_over_font(
    input  wire        clk,
    input  wire [15:0] addr,            
    output reg  [63:0]  char_line_pixels 
);

    // signal declaration
    reg [63:0] data;

// body
always @(posedge clk)
    char_line_pixels <= data;

always @* begin
    case (addr)
        //code x00
        16'h0000: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0001: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0002: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0003: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0004: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0005: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0006: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0007: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0008: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0009: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h000f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0010: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0011: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0012: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0013: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0014: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0015: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0016: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0017: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0018: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0019: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h001f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0020: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0021: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0022: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0023: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0024: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0025: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0026: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0027: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
       
        16'h0028: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0029: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h002f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0030: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0031: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0032: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0033: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0034: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0035: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0036: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0037: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h0038: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h0039: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h003f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x41
        16'h4100: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4101: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4102: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4103: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4104: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4105: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4106: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
        16'h4107: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;
       
        16'h4108: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000;
        16'h4109: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000;
        16'h410a: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000;
        16'h410b: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000; 
        16'h410c: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000; 
        16'h410d: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000; 
        16'h410e: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000; 
        16'h410f: data = 64'b00000000_11111111_11111111_00000000_11111111_11111111_00000000_00000000; 
       
        16'h4110: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4111: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4112: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4113: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4114: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4115: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4116: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4117: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
       
        16'h4118: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4119: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h411f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
       
        16'h4120: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4121: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4122: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4123: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4124: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4125: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4126: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4127: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        
        16'h4128: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4129: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h412f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
       
        16'h4130: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h4131: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;  
        16'h4132: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4133: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4134: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4135: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4136: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4137: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
       
        16'h4138: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4139: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h413f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
       
        //code x45
        16'h4500: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4501: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4502: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4503: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4504: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4505: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4506: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4507: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        
        16'h4508: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4509: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h450a: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h450b: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h450c: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h450d: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h450e: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h450f: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        
        16'h4510: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4511: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4512: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4513: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4514: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4515: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4516: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4517: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h4518: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h4519: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451a: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451b: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451c: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451d: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451e: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h451f: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000;
        
        16'h4520: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4521: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4522: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4523: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4524: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4525: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4526: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4527: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        
        16'h4528: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4529: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;  
        16'h452a: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h452b: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h452c: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h452d: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;  
        16'h452e: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h452f: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000;  
        
        16'h4530: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4531: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4532: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4533: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4534: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4535: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4536: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4537: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        
        16'h4538: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h4539: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h453a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h453b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h453c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h453d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h453e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h453f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        
        //code x47
        16'h4700: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4701: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4702: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4703: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4704: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4705: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4706: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4707: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h4708: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h4709: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470a: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470b: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470c: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470d: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470e: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        16'h470f: data = 64'b00000000_11111111_11111111_00000000_00000000_00000000_00000000_00000000; 
        
        16'h4710: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4711: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4712: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4713: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4714: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4715: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4716: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4717: data = 64'b11111111_11111111_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        16'h4718: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h4719: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471a: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471b: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471c: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471d: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471e: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h471f: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 

        16'h4720: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4721: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4722: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4723: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4724: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4725: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4726: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4727: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4728: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h4729: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472a: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472b: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472c: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472d: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472e: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 
        16'h472f: data = 64'b00000000_11111111_11111111_00000000_00000000_11111111_11111111_00000000; 

        16'h4730: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4731: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4732: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4733: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4734: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4735: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4736: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4737: data = 64'b00000000_00000000_11111111_11111111_11111111_11111111_11111111_00000000; 

        16'h4738: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4739: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h473f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 

        //code x4D
        16'h4d00: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d01: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d02: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d03: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d04: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d05: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d06: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h4d07: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;

        16'h4d08: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d09: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d0a: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000; 
        16'h4d0b: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d0c: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d0d: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d0e: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;
        16'h4d0f: data = 64'b11111111_11111111_11111111_00000000_11111111_11111111_11111111_00000000;

        16'h4d10: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d11: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d12: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d13: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;        
        16'h4d14: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d15: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d16: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d17: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        
        16'h4d18: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d19: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d1a: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d1b: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d1c: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d1d: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000; 
        16'h4d1e: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        16'h4d1f: data = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_00000000;
        
        16'h4d20: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d21: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d22: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d23: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d24: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d25: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d26: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        16'h4d27: data = 64'b11111111_11111111_00000000_11111111_00000000_11111111_11111111_00000000;
        
        16'h4d28: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d29: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d2f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4d30: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d31: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d32: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d33: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d34: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d35: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d36: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4d37: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        
        16'h4d38: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d39: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4d3f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        
        //code x4F
        16'h4f00: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f01: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f02: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f03: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f04: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f05: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f06: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f07: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h4f08: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f09: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f0f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f10: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f11: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f12: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f13: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f14: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f15: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f16: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f17: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f18: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f19: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f1f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f20: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f21: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f22: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f23: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f24: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f25: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f26: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f27: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f28: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f29: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h4f2f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h4f30: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f31: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f32: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f33: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f34: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f35: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f36: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h4f37: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h4f38: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f39: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h4f3f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        //code x52
        16'h5200: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5201: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5202: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5203: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5204: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5205: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5206: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5207: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h5208: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5209: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h520a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h520b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h520c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h520d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h520e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h520f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        
        16'h5210: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5211: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5212: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5213: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5214: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5215: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5216: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5217: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        
        16'h5218: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;
        16'h5219: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;
        16'h521a: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h521b: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h521c: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;
        16'h521d: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000;
        16'h521e: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        16'h521f: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_11111111_00000000; 
        
        16'h5220: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5221: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5222: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5223: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5224: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5225: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5226: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5227: data = 64'b11111111_11111111_11111111_11111111_11111111_00000000_00000000_00000000; 
        
        16'h5228: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000; 
        16'h5229: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000;   
        16'h522a: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000; 
        16'h522b: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000; 
        16'h522c: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000; 
        16'h522d: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000;  
        16'h522e: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000; 
        16'h522f: data = 64'b11111111_11111111_00000000_00000000_11111111_11111111_00000000_00000000;   
        
        16'h5230: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5231: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5232: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5233: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5234: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5235: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5236: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5237: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        
        16'h5238: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h5239: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h523a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h523b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h523c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h523d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h523e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h523f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        
        //code x56
        16'h5600: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5601: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5602: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5603: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5604: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5605: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5606: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5607: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5608: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000;
        16'h5609: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h560f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5610: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5611: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5612: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5613: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5614: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5615: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5616: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5617: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5618: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h5619: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561a: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561b: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561c: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561d: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561e: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        16'h561f: data = 64'b11111111_11111111_00000000_00000000_00000000_11111111_11111111_00000000; 
        
        16'h5620: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5621: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5622: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5623: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5624: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5625: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5626: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        16'h5627: data = 64'b00000000_11111111_11111111_11111111_11111111_11111111_00000000_00000000; 
        
        16'h5628: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h5629: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;  
        16'h562a: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h562b: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h562c: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h562d: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000;  
        16'h562e: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        16'h562f: data = 64'b00000000_00000000_11111111_11111111_11111111_00000000_00000000_00000000; 
        
        16'h5630: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        16'h5631: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        16'h5632: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        16'h5633: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000;
        16'h5634: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        16'h5635: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000;
        16'h5636: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        16'h5637: data = 64'b00000000_00000000_00000000_11111111_00000000_00000000_00000000_00000000; 
        
        16'h5638: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h5639: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h563a: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h563b: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
        16'h563c: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h563d: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h563e: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        16'h563f: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; 
        
        default: data = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
    endcase
end

endmodule
