`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_small_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arcade_small_font(
        input  wire        clk,
        input  wire [15:0] addr,            
        output reg  [39:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [39:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
        //code x00
16'h0000: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0001: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0002: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0003: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0004: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
                 
16'h0005: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0006: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0007: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0008: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0009: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                
16'h000a: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h000b: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h000c: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h000d: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h000e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h000f: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0010: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0011: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0012: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0013: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h0014: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0015: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0016: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0017: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0018: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;

16'h0019: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h001a: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h001b: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h001c: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h001d: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h001e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h001f: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0020: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0021: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0022: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h0023: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0024: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0025: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0026: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h0027: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
                
                
                
    //code x3A
16'h3a00: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a01: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a02: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a03: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a04: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
       
16'h3a05: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a06: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a07: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a08: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a09: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        
16'h3a0a: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a0b: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a0c: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a0d: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a0e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h3a0f: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a10: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a11: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a12: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a13: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 

16'h3a14: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a15: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a16: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a17: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a18: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;

16'h3a19: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a1a: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a1b: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a1c: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 
16'h3a1d: data = 40'b00000_11111_00000_00000_00000_00000_00000_00000; 

16'h3a1e: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a1f: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a20: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a21: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a22: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

16'h3a23: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a24: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a25: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a26: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h3a27: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;
               
                
                
                
                
                
                       //code x41
16'h4100: data = 40'b00000_00000_11111_11111_11111_00000_00000_00000;
16'h4101: data = 40'b00000_00000_11111_11111_11111_00000_00000_00000;
16'h4102: data = 40'b00000_00000_11111_11111_11111_00000_00000_00000;
16'h4103: data = 40'b00000_00000_11111_11111_11111_00000_00000_00000;
16'h4104: data = 40'b00000_00000_11111_11111_11111_00000_00000_00000;

16'h4105: data = 40'b00000_11111_11111_00000_11111_11111_00000_00000;
16'h4106: data = 40'b00000_11111_11111_00000_11111_11111_00000_00000; 
16'h4107: data = 40'b00000_11111_11111_00000_11111_11111_00000_00000;
16'h4108: data = 40'b00000_11111_11111_00000_11111_11111_00000_00000;
16'h4109: data = 40'b00000_11111_11111_00000_11111_11111_00000_00000;

16'h410a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h410b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h410c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h410d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h410e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h410f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4110: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4111: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4112: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4113: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4114: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4115: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4116: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000; 
16'h4117: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;  
16'h4118: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000; 

16'h4119: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h411a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h411b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h411c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h411d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h411e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h411f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4120: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4121: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4122: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4123: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4124: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4125: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4126: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4127: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

       
       
       
                                    //code x43
16'h4300: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h4301: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
16'h4302: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
16'h4303: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
16'h4304: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;

16'h4305: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h4306: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h4307: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h4308: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h4309: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;

16'h430a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h430b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h430c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h430d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h430e: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;

16'h430f: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h4310: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4311: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h4312: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4313: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 

16'h4314: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4315: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4316: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4317: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4318: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 

16'h4319: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h431a: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h431b: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h431c: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h431d: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 

16'h431e: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h431f: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h4320: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h4321: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h4322: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;

16'h4323: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4324: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4325: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4326: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4327: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

                
                
                
                
                
                
                          //code x45
16'h4500: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4501: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4502: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4503: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4504: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;

16'h4505: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4506: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4507: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4508: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4509: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  

16'h450a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h450b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h450c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h450d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h450e: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  

16'h450f: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h4510: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h4511: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h4512: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h4513: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 

16'h4514: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4515: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4516: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h4517: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;   
16'h4518: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 

16'h4519: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h451a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h451b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h451c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h451d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 

16'h451e: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h451f: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4520: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4521: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;
16'h4522: data = 40'b11111_11111_11111_11111_11111_11111_11111_00000;

16'h4523: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4524: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4525: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4526: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4527: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
                 
                        //code x4F
16'h4f00: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f01: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f02: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f03: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f04: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h4f05: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f06: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f07: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f08: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f09: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4f0a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f0b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f0c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f0d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f0e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4f0f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f10: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f11: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f12: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f13: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4f14: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f15: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f16: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f17: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;   
16'h4f18: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4f19: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f1a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f1b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f1c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h4f1d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h4f1e: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h4f1f: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f20: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f21: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h4f22: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h4f23: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4f24: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4f25: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4f26: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h4f27: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 

  
  
  
                          //code x50
16'h5000: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5001: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5002: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5003: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5004: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;

16'h5005: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5006: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5007: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5008: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5009: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;

16'h500a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h500b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h500c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h500d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h500e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;

16'h500f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5010: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5011: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5012: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5013: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;

16'h5014: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5015: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5016: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;
16'h5017: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000; 
16'h5018: data = 40'b11111_11111_11111_11111_11111_11111_00000_00000;  

16'h5019: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h501a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h501b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;   
16'h501c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h501d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  

16'h501e: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h501f: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h5020: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h5021: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;  
16'h5022: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 

16'h5023: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5024: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5025: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5026: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5027: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 





         
                          //code x52
16'h5200: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5201: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5202: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5203: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5204: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h5205: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5206: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5207: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5208: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5209: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;  

16'h520a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;  
16'h520b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h520c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h520d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h520e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;  

16'h520f: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
16'h5210: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 
16'h5211: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000;  
16'h5212: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000;  
16'h5213: data = 40'b11111_11111_00000_00000_11111_11111_11111_00000; 

16'h5214: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h5215: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h5216: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 
16'h5217: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000;   
16'h5218: data = 40'b11111_11111_11111_11111_11111_00000_00000_00000; 

16'h5219: data = 40'b11111_11111_00000_00000_11111_11111_00000_00000; 
16'h521a: data = 40'b11111_11111_00000_00000_11111_11111_00000_00000; 
16'h521b: data = 40'b11111_11111_00000_00000_11111_11111_00000_00000; 
16'h521c: data = 40'b11111_11111_00000_00000_11111_11111_00000_00000; 
16'h521d: data = 40'b11111_11111_00000_00000_11111_11111_00000_00000; 

16'h521e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h521f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5220: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5221: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;
16'h5222: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;

16'h5223: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5224: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5225: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5226: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5227: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;




         
    //code x53
16'h5300: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h5301: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;  
16'h5302: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;  
16'h5303: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;  
16'h5304: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h5305: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5306: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5307: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5308: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5309: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h530a: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h530b: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h530c: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h530d: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000; 
16'h530e: data = 40'b11111_11111_00000_00000_00000_00000_00000_00000;

16'h530f: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;  
16'h5310: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5311: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h5312: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5313: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h5314: data = 40'b00000_00000_00000_00000_00000_11111_11111_00000; 
16'h5315: data = 40'b00000_00000_00000_00000_00000_11111_11111_00000; 
16'h5316: data = 40'b00000_00000_00000_00000_00000_11111_11111_00000; 
16'h5317: data = 40'b00000_00000_00000_00000_00000_11111_11111_00000;  
16'h5318: data = 40'b00000_00000_00000_00000_00000_11111_11111_00000; 

16'h5319: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;  
16'h531a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h531b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h531c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h531d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h531e: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h531f: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h5320: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h5321: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h5322: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h5323: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5324: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5325: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5326: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5327: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;   


        
        
        
        
        
        
        //code x54
16'h5400: data = 40'b00000_11111_11111_11111_11111_11111_11111_00000;
16'h5401: data = 40'b00000_11111_11111_11111_11111_11111_11111_00000; 
16'h5402: data = 40'b00000_11111_11111_11111_11111_11111_11111_00000; 
16'h5403: data = 40'b00000_11111_11111_11111_11111_11111_11111_00000;
16'h5404: data = 40'b00000_11111_11111_11111_11111_11111_11111_00000;
  
16'h5405: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5406: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5407: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5408: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5409: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 

16'h540a: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h540b: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h540c: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h540d: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h540e: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
 
16'h540f: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5410: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5411: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5412: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5413: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 

16'h5414: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5415: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5416: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5417: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5418: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  

16'h5419: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h541a: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h541b: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h541c: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h541d: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  

16'h541e: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h541f: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5420: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5421: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5422: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;
 
16'h5423: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5424: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5425: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5426: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5427: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        


         
         
        
                                  //code x55
16'h5500: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5501: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5502: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5503: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5504: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h5505: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5506: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5507: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5508: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5509: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h550a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h550b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h550c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h550d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h550e: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h550f: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5510: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5511: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5512: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5513: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h5514: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5515: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5516: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h5517: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000;   
16'h5518: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h5519: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h551a: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h551b: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h551c: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 
16'h551d: data = 40'b11111_11111_00000_00000_00000_11111_11111_00000; 

16'h551e: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000; 
16'h551f: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5520: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5521: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;
16'h5522: data = 40'b00000_11111_11111_11111_11111_11111_00000_00000;

16'h5523: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5524: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5525: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5526: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5527: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 








  //code x59
16'h5900: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h5901: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h5902: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000; 
16'h5903: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h5904: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
  
16'h5905: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h5906: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h5907: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;  
16'h5908: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h5909: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;

16'h590a: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h590b: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h590c: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h590d: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
16'h590e: data = 40'b00000_11111_11111_00000_00000_11111_11111_00000;
 
16'h590f: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h5910: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;   
16'h5911: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 
16'h5912: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000;  
16'h5913: data = 40'b00000_00000_11111_11111_11111_11111_00000_00000; 

16'h5914: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5915: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h5916: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5917: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5918: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  

16'h5919: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h591a: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h591b: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  
16'h591c: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h591d: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;  

16'h591e: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h591f: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5920: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5921: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000; 
16'h5922: data = 40'b00000_00000_00000_11111_11111_00000_00000_00000;
 
16'h5923: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5924: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5925: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5926: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
16'h5927: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000; 
        
 default: data = 40'b00000_00000_00000_00000_00000_00000_00000_00000;

        endcase

endmodule

