`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_numbers_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Ma�a czcionka dla cyfr
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// Wzorowano na czcionce Arcade Classic
//////////////////////////////////////////////////////////////////////////////////


module arcade_numbers_font(
    input  wire        clk,
    input  wire [15:0] addr,            
    output reg  [31:0] char_line_pixels 
);
    
    // signal declaration
    reg [31:0] data;

// body
always @(posedge clk)
    char_line_pixels <= data;

always @* begin
    case (addr)
        //code x00
        16'h0000: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0001: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0002: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0003: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
             
        16'h0004: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;      
        16'h0005: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h0006: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h0007: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
                 
        16'h0008: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h0009: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h000a: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h000b: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
               
        16'h000c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h000d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h000e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;     
        16'h000f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
               
        16'h0010: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h0011: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0012: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0013: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
                       
        16'h0014: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h0015: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0016: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h0017: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
               
        16'h0018: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;   
        16'h0019: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h001a: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h001b: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
               
        16'h001c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h001d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;      
        16'h001e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h001f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 

        //code x30
        16'h3000: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3001: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3002: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3003: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        
        16'h3004: data = 32'b0000_1111_0000_0000_1111_1111_0000_0000;
        16'h3005: data = 32'b0000_1111_0000_0000_1111_1111_0000_0000; 
        16'h3006: data = 32'b0000_1111_0000_0000_1111_1111_0000_0000;
        16'h3007: data = 32'b0000_1111_0000_0000_1111_1111_0000_0000; 
        
        16'h3008: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3009: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h300a: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h300b: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h300c: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h300d: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h300e: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h300f: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h3010: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3011: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3012: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3013: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h3014: data = 32'b0000_1111_1111_0000_0000_1111_0000_0000; 
        16'h3015: data = 32'b0000_1111_1111_0000_0000_1111_0000_0000; 
        16'h3016: data = 32'b0000_1111_1111_0000_0000_1111_0000_0000; 
        16'h3017: data = 32'b0000_1111_1111_0000_0000_1111_0000_0000;   
        
        16'h3018: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000; 
        16'h3019: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000; 
        16'h301a: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000; 
        16'h301b: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000; 
        
        16'h301c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h301d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h301e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h301f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        
        //code x31
        16'h3100: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3101: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3102: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3103: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h3104: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3105: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3106: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000;
        16'h3107: data = 32'b0000_0000_1111_1111_1111_0000_0000_0000; 
        
        16'h3108: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3109: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h310a: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h310b: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h310c: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h310d: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h310e: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h310f: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h3110: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;  
        16'h3111: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3112: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3113: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h3114: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000; 
        16'h3115: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;  
        16'h3116: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000; 
        16'h3117: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000; 
        
        16'h3118: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        16'h3119: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        16'h311a: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        16'h311b: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        
        16'h311c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h311d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;  
        16'h311e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h311f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        
        //code x32
        16'h3200: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;
        16'h3201: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;
        16'h3202: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;
        16'h3203: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;
        
        16'h3204: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3205: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3206: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3207: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        
        16'h3208: data = 32'b0000_0000_0000_00000_1111_1111_1111_0000;
        16'h3209: data = 32'b0000_0000_0000_00000_1111_1111_1111_0000;
        16'h320a: data = 32'b0000_0000_0000_00000_1111_1111_1111_0000; 
        16'h320b: data = 32'b0000_0000_0000_00000_1111_1111_1111_0000; 
        
        16'h320c: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000; 
        16'h320d: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;  
        16'h320e: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000; 
        16'h320f: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000; 
        
        16'h3210: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        16'h3211: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;   
        16'h3212: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        16'h3213: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        
        16'h3214: data = 32'b1111_1111_1111_0000_0000_0000_0000_0000; 
        16'h3215: data = 32'b1111_1111_1111_0000_0000_0000_0000_0000; 
        16'h3216: data = 32'b1111_1111_1111_0000_0000_0000_0000_0000; 
        16'h3217: data = 32'b1111_1111_1111_0000_0000_0000_0000_0000; 
        
        16'h3218: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h3219: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h321a: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h321b: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;  
        
        16'h321c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h321d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h321e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h321f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        
        //code x33
        16'h3300: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;
        16'h3301: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;
        16'h3302: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;
        16'h3303: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        
        16'h3304: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3305: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3306: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3307: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        
        16'h3308: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h3309: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h330a: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h330b: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h330c: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h330d: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h330e: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h330f: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000; 
        
        16'h3310: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        16'h3311: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        16'h3312: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        16'h3313: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        
        16'h3314: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3315: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3316: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3317: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h3318: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h3319: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h331a: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h331b: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        
        16'h331c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h331d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h331e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h331f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        
        //code x34
        16'h3400: data = 32'b0000_0000_0000_1111_1111_1111_0000_0000;
        16'h3401: data = 32'b0000_0000_0000_1111_1111_1111_0000_0000;
        16'h3402: data = 32'b0000_0000_0000_1111_1111_1111_0000_0000;
        16'h3403: data = 32'b0000_0000_0000_1111_1111_1111_0000_0000;
        
        16'h3404: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3405: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3406: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3407: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        
        16'h3408: data = 32'b0000_1111_1111_0000_1111_1111_0000_0000;
        16'h3409: data = 32'b0000_1111_1111_0000_1111_1111_0000_0000;
        16'h340a: data = 32'b0000_1111_1111_0000_1111_1111_0000_0000;  
        16'h340b: data = 32'b0000_1111_1111_0000_1111_1111_0000_0000; 
        
        16'h340c: data = 32'b1111_1111_0000_0000_1111_1111_0000_0000;  
        16'h340d: data = 32'b1111_1111_0000_0000_1111_1111_0000_0000; 
        16'h340e: data = 32'b1111_1111_0000_0000_1111_1111_0000_0000; 
        16'h340f: data = 32'b1111_1111_0000_0000_1111_1111_0000_0000; 
        
        16'h3410: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h3411: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h3412: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        16'h3413: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000; 
        
        16'h3414: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3415: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3416: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3417: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;  
        
        16'h3418: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h3419: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h341a: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h341b: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        
        16'h341c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h341d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h341e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h341f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        
        //code x35
        16'h3500: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3501: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3502: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3503: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        
        16'h3504: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000;
        16'h3505: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000;
        16'h3506: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000;
        16'h3507: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000;
        
        16'h3508: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000;
        16'h3509: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000;
        16'h350a: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000;
        16'h350b: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000;
        
        16'h350c: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        16'h350d: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        16'h350e: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        16'h350f: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        
        16'h3510: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        16'h3511: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;  
        16'h3512: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;  
        16'h3513: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;  
        
        16'h3514: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;  
        16'h3515: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;  
        16'h3516: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;  
        16'h3517: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;   
        
        16'h3518: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;  
        16'h3519: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h351a: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h351b: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        
        16'h351c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h351d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h351e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h351f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
       
        //code x36
        16'h3600: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3601: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3602: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        16'h3603: data = 32'b0000_0000_1111_1111_1111_1111_0000_0000;
        
        16'h3604: data = 32'b0000_1111_1111_0000_0000_0000_0000_0000;
        16'h3605: data = 32'b0000_1111_1111_0000_0000_0000_0000_0000; 
        16'h3606: data = 32'b0000_1111_1111_0000_0000_0000_0000_0000; 
        16'h3607: data = 32'b0000_1111_1111_0000_0000_0000_0000_0000; 
        
        16'h3608: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000; 
        16'h3609: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000; 
        16'h360a: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000; 
        16'h360b: data = 32'b1111_1111_0000_0000_0000_0000_0000_0000; 
        
        16'h360c: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000; 
        16'h360d: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000; 
        16'h360e: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000; 
        16'h360f: data = 32'b1111_1111_1111_1111_1111_1111_0000_0000;
        
        16'h3610: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3611: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3612: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3613: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        
        16'h3614: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3615: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3616: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3617: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;   
        
        16'h3618: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h3619: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h361a: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h361b: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        
        16'h361c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h361d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h361e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h361f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        
        //code x37
        16'h3700: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3701: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3702: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        16'h3703: data = 32'b1111_1111_1111_1111_1111_1111_1111_0000;
        
        16'h3704: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3705: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3706: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3707: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h3708: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h3709: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h370a: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        16'h370b: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;
        
        16'h370c: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h370d: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h370e: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        16'h370f: data = 32'b0000_0000_0000_1111_1111_0000_0000_0000;
        
        16'h3710: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3711: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3712: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3713: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        
        16'h3714: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3715: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3716: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3717: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        
        16'h3718: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h3719: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h371a: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000;
        16'h371b: data = 32'b0000_0000_1111_1111_0000_0000_0000_0000; 
        
        16'h371c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h371d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h371e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h371f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        
        //code x38
        16'h3800: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;
        16'h3801: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;
        16'h3802: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;
        16'h3803: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;
        
        16'h3804: data = 32'b1111_1111_0000_0000_0000_1111_0000_0000;
        16'h3805: data = 32'b1111_1111_0000_0000_0000_1111_0000_0000; 
        16'h3806: data = 32'b1111_1111_0000_0000_0000_1111_0000_0000; 
        16'h3807: data = 32'b1111_1111_0000_0000_0000_1111_0000_0000; 
        
        16'h3808: data = 32'b1111_1111_1111_0000_0000_1111_0000_0000; 
        16'h3809: data = 32'b1111_1111_1111_0000_0000_1111_0000_0000;  
        16'h380a: data = 32'b1111_1111_1111_0000_0000_1111_0000_0000;  
        16'h380b: data = 32'b1111_1111_1111_0000_0000_1111_0000_0000;  
        
        16'h380c: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;  
        16'h380d: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;  
        16'h380e: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;  
        16'h380f: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000;
        
        16'h3810: data = 32'b1111_0000_0000_1111_1111_1111_1111_0000;
        16'h3811: data = 32'b1111_0000_0000_1111_1111_1111_1111_0000; 
        16'h3812: data = 32'b1111_0000_0000_1111_1111_1111_1111_0000;
        16'h3813: data = 32'b1111_0000_0000_1111_1111_1111_1111_0000;
        
        16'h3814: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3815: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3816: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3817: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;  
        
        16'h3818: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h3819: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h381a: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h381b: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        
        16'h381c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h381d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h381e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        16'h381f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        
        //code x39
        16'h3900: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000; 
        16'h3901: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;  
        16'h3902: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;  
        16'h3903: data = 32'b0000_1111_1111_1111_1111_1111_0000_0000;  
        
        16'h3904: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        16'h3905: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3906: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3907: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        
        16'h3908: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h3909: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h390a: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000; 
        16'h390b: data = 32'b1111_1111_0000_0000_0000_1111_1111_0000;
        
        16'h390c: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000; 
        16'h390d: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000; 
        16'h390e: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;
        16'h390f: data = 32'b0000_1111_1111_1111_1111_1111_1111_0000;  
        
        16'h3910: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        16'h3911: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000; 
        16'h3912: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        16'h3913: data = 32'b0000_0000_0000_0000_0000_1111_1111_0000;
        
        16'h3914: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h3915: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h3916: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000; 
        16'h3917: data = 32'b0000_0000_0000_0000_1111_1111_0000_0000;  
        
        16'h3918: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        16'h3919: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        16'h391a: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        16'h391b: data = 32'b0000_1111_1111_1111_1111_0000_0000_0000; 
        
        16'h391c: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h391d: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h391e: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        16'h391f: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
        
        default: data = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    endcase
end

endmodule
