`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.07.2022 18:45:55
// Design Name: 
// Module Name: arcade_big_font
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arcade_you_win_font(
        input  wire        clk,
        input  wire [15:0] addr,            
        output reg  [79:0]  char_line_pixels 
    );

    // signal declaration
    reg [79:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
        //code x00
                16'h0000: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0001: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0002: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0003: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0004: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0005: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0006: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0007: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0008: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0009: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h000a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h000f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0010: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0011: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0012: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0013: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
              
                16'h0014: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0015: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0016: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0017: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0018: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0019: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
       
                16'h001e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h001f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0020: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0021: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0022: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0023: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0024: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0025: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0026: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0027: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h0028: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0029: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h002f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0030: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0031: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        
                16'h0032: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0033: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0034: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0035: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0036: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0037: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0038: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0039: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                
                16'h003c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h003f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0040: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0041: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0042: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0043: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0044: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0045: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                
                16'h0046: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0047: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0048: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h0049: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h004f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;

//code x4F
     16'h4f00: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f01: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f02: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f03: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f04: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f05: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f06: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f07: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f08: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f09: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     
     16'h4f0a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f0f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f10: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f11: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f12: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f13: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
    
     16'h4f14: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f15: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f16: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f17: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f18: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f19: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     
     16'h4f1e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f1f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f20: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f21: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f22: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f23: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f24: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f25: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f26: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f27: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     
     16'h4f28: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f29: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f2f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f30: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f31: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 

     16'h4f32: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f33: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f34: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f35: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f36: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f37: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f38: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f39: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f3a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
     16'h4f3b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
    
     16'h4f3c: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3d: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3e: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f3f: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f40: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f41: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f42: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f43: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f44: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     16'h4f45: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
     
     16'h4f46: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f47: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f48: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f49: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
     16'h4f4f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;


           //code x49
                            16'h4900: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4901: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4902: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                            16'h4903: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4904: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4905: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4906: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4907: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4908: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4909: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                            
                            16'h490a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h490b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h490c: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;   
                            16'h490d: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h490e: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h490f: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4910: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4911: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4912: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4913: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            
                            16'h4914: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4915: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4916: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;   
                            16'h4917: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4918: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4919: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h491a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h491b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h491c: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h491d: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            
                            16'h491e: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h491f: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4920: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;   
                            16'h4921: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4922: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4923: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4924: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4925: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4926: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4927: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;
                          
                            16'h4928: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4929: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
                            16'h492a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
                            16'h492b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h492c: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h492d: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h492e: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h492f: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4930: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4931: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;
                                     
                            16'h4932: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4933: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4934: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;   
                            16'h4935: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4936: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4937: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4938: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h4939: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h493a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                            16'h493b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
                              
                            16'h493c: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h493d: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h493e: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                            16'h493f: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4940: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4941: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4942: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4943: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4944: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                            16'h4945: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                                     
                            16'h4946: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h4947: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h4948: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h4949: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                            16'h494f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
      //code x4e
                                       16'h4e00: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e01: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                                       16'h4e02: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                                       16'h4e03: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                                       16'h4e04: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e05: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e06: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e07: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e08: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                                       16'h4e09: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                     
                                       16'h4e0a: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e0b: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e0c: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e0d: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e0e: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e0f: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e10: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e11: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e12: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e13: data = 80'b1111111111_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                      
                                       16'h4e14: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e15: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e16: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e17: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e18: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e19: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e1a: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e1b: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e1c: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e1d: data = 80'b1111111111_1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_0000000000; 
                                       
                                       16'h4e1e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e1f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e20: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e21: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e22: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e23: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e24: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e25: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e26: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e27: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       
                                       16'h4e28: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;  
                                       16'h4e29: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;   
                                       16'h4e2a: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;  
                                       16'h4e2b: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;  
                                       16'h4e2c: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e2d: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;   
                                       16'h4e2e: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e2f: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e30: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e31: data = 80'b1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000;  
                                  
                                       16'h4e32: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e33: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                       16'h4e34: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                       16'h4e35: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                       16'h4e36: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e37: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e38: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                       16'h4e39: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000; 
                                       16'h4e3a: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                       16'h4e3b: data = 80'b1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_1111111111_0000000000;
                                      
                                       16'h4e3c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e3d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e3e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e3f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e40: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e41: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e42: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e43: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e44: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                                       16'h4e45: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;  
                                  
                                       16'h4e46: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e47: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e48: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e49: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                                       16'h4e4f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                             
              
              
                       //code x55
                         16'h5500: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5501: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                         16'h5502: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5503: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                         16'h5504: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5505: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5506: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5507: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5508: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5509: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         
                         16'h550a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h550b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h550c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h550d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h550e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h550f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5510: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5511: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5512: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5513: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                        
                         16'h5514: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5515: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5516: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5517: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5518: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5519: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h551a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h551b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h551c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h551d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         
                         16'h551e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h551f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5520: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5521: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5522: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5523: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5524: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5525: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5526: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5527: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         
                         16'h5528: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5529: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h552f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5530: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5531: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                     
                         16'h5532: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5533: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5534: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5535: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5536: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5537: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5538: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h5539: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h553a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                         16'h553b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                        
                         16'h553c: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h553d: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h553e: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h553f: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5540: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5541: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5542: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5543: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5544: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         16'h5545: data = 80'b0000000000_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
                         
                         16'h5546: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h5547: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h5548: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h5549: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                         16'h554f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
   
//code x57
                16'h5700: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5701: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                16'h5702: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                16'h5703: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                16'h5704: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5705: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5706: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5707: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5708: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;
                16'h5709: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
              
                16'h570a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h570b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h570c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h570d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h570e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h570f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5710: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5711: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5712: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5713: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
               
                16'h5714: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5715: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5716: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5717: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5718: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5719: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h571a: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h571b: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h571c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h571d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                
                16'h571e: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h571f: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5720: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5721: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5722: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5723: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5724: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5725: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5726: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                16'h5727: data = 80'b1111111111_1111111111_0000000000_1111111111_0000000000_1111111111_1111111111_0000000000; 
                
                16'h5728: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                16'h5729: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;   
                16'h572a: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                16'h572b: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
                16'h572c: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                16'h572d: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;   
                16'h572e: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                16'h572f: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                16'h5730: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000; 
                16'h5731: data = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_0000000000;  
           
                16'h5732: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000; 
                16'h5733: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                16'h5734: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                16'h5735: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                16'h5736: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000; 
                16'h5737: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000; 
                16'h5738: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                16'h5739: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000; 
                16'h573a: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                16'h573b: data = 80'b1111111111_1111111111_1111111111_0000000000_1111111111_1111111111_1111111111_0000000000;
                
                16'h573c: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h573d: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h573e: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h573f: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5740: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5741: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5742: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5743: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5744: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000; 
                16'h5745: data = 80'b1111111111_1111111111_0000000000_0000000000_0000000000_1111111111_1111111111_0000000000;  
                
                16'h5746: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h5747: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h5748: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h5749: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
                16'h574f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;


                    //code x59
        16'h5900: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5901: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000;  
        16'h5902: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5903: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5904: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5905: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5906: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5907: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5908: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5909: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        
        16'h590a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h590b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h590c: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h590d: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h590e: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h590f: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5910: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5911: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5912: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5913: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
       
        16'h5914: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5915: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5916: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5917: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5918: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h5919: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h591a: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h591b: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 
        16'h591c: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000;  
        16'h591d: data = 80'b0000000000_1111111111_1111111111_0000000000_0000000000_1111111111_1111111111_0000000000; 

        16'h591e: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h591f: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000;  
        16'h5920: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000;  
        16'h5921: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5922: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5923: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5924: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5925: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5926: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        16'h5927: data = 80'b0000000000_0000000000_1111111111_1111111111_1111111111_1111111111_0000000000_0000000000; 
        
        16'h5928: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5929: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h592a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
        16'h592b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h592c: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h592d: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h592e: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h592f: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5930: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5931: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;
        
        16'h5932: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5933: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5934: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
        16'h5935: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5936: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5937: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5938: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5939: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h593a: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h593b: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 

        16'h593c: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h593d: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h593e: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
        16'h593f: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5940: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5941: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5942: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5943: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5944: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000; 
        16'h5945: data = 80'b0000000000_0000000000_0000000000_1111111111_1111111111_0000000000_0000000000_0000000000;  
       
        16'h5946: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h5947: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h5948: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h5949: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594a: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594b: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594c: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594d: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594e: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000; 
        16'h594f: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;

 	default: data = 80'b0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000;
        endcase

endmodule
